-- Copyright 2018 Jonas Fuhrmann. All rights reserved.
--
-- This project is dual licensed under GNU General Public License version 3
-- and a commercial license available on request.
---------------------------------------------------------------------------
-- For non commercial use only:
-- This file is part of tinyTPU.
-- 
-- tinyTPU is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
-- 
-- tinyTPU is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with tinyTPU. If not, see <http://www.gnu.org/licenses/>.

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

PACKAGE TPU_PACK IS
    CONSTANT BYTE_WIDTH : NATURAL := 8;
    CONSTANT EXTENDED_BYTE_WIDTH : NATURAL := BYTE_WIDTH + 1;

    SUBTYPE BYTE_TYPE IS STD_LOGIC_VECTOR(BYTE_WIDTH - 1 DOWNTO 0);
    SUBTYPE EXTENDED_BYTE_TYPE IS STD_LOGIC_VECTOR(EXTENDED_BYTE_WIDTH - 1 DOWNTO 0);
    SUBTYPE MUL_HALFWORD_TYPE IS STD_LOGIC_VECTOR(2 * EXTENDED_BYTE_WIDTH - 1 DOWNTO 0);
    SUBTYPE HALFWORD_TYPE IS STD_LOGIC_VECTOR(2 * BYTE_WIDTH - 1 DOWNTO 0);
    SUBTYPE WORD_TYPE IS STD_LOGIC_VECTOR(4 * BYTE_WIDTH - 1 DOWNTO 0);

    TYPE INTEGER_ARRAY_TYPE IS ARRAY(INTEGER RANGE <>) OF INTEGER;
    TYPE BIT_ARRAY_2D_TYPE IS ARRAY(NATURAL RANGE <>, NATURAL RANGE <>) OF STD_LOGIC;
    TYPE BYTE_ARRAY_TYPE IS ARRAY(NATURAL RANGE <>) OF BYTE_TYPE;
    TYPE BYTE_ARRAY_2D_TYPE IS ARRAY(NATURAL RANGE <>, NATURAL RANGE <>) OF BYTE_TYPE;
    TYPE EXTENDED_BYTE_ARRAY IS ARRAY(NATURAL RANGE <>) OF EXTENDED_BYTE_TYPE;
    TYPE HALFWORD_ARRAY_TYPE IS ARRAY(NATURAL RANGE <>) OF HALFWORD_TYPE;
    TYPE WORD_ARRAY_TYPE IS ARRAY(NATURAL RANGE <>) OF WORD_TYPE;
    TYPE WORD_ARRAY_2D_TYPE IS ARRAY(NATURAL RANGE <>, NATURAL RANGE <>) OF WORD_TYPE;

    -- Good for readable testbenches
    TYPE INTEGER_ARRAY_2D_TYPE IS ARRAY(NATURAL RANGE <>, NATURAL RANGE <>) OF INTEGER;

    -- Type for activation
    SUBTYPE ACTIVATION_BIT_TYPE IS STD_LOGIC_VECTOR(3 DOWNTO 0);
    TYPE ACTIVATION_TYPE IS (NO_ACTIVATION, RELU, RELU6, CRELU, ELU, SELU, SOFTPLUS, SOFTSIGN, DROPOUT, SIGMOID, TANH);
    -- Conversion functions
    FUNCTION BITS_TO_ACTIVATION(BITVECTOR : ACTIVATION_BIT_TYPE) RETURN ACTIVATION_TYPE;
    FUNCTION ACTIVATION_TO_BITS(ACTIVATION_FUNCTION : ACTIVATION_TYPE) RETURN ACTIVATION_BIT_TYPE;

    FUNCTION BITS_TO_BYTE_ARRAY(BITVECTOR : STD_LOGIC_VECTOR) RETURN BYTE_ARRAY_TYPE;
    FUNCTION BYTE_ARRAY_TO_BITS(BYTE_ARRAY : BYTE_ARRAY_TYPE) RETURN STD_LOGIC_VECTOR;

    FUNCTION BITS_TO_WORD_ARRAY(BITVECTOR : STD_LOGIC_VECTOR) RETURN WORD_ARRAY_TYPE;
    FUNCTION WORD_ARRAY_TO_BITS(WORD_ARRAY : WORD_ARRAY_TYPE) RETURN STD_LOGIC_VECTOR;

    -- Control types
    CONSTANT BUFFER_ADDRESS_WIDTH : NATURAL := 24;
    CONSTANT ACCUMULATOR_ADDRESS_WIDTH : NATURAL := 16;
    CONSTANT WEIGHT_ADDRESS_WIDTH : NATURAL := BUFFER_ADDRESS_WIDTH + ACCUMULATOR_ADDRESS_WIDTH;
    CONSTANT LENGTH_WIDTH : NATURAL := 32;
    CONSTANT OP_CODE_WIDTH : NATURAL := 8;
    CONSTANT INSTRUCTION_WIDTH : NATURAL := WEIGHT_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH;

    SUBTYPE BUFFER_ADDRESS_TYPE IS STD_LOGIC_VECTOR(BUFFER_ADDRESS_WIDTH - 1 DOWNTO 0);
    SUBTYPE ACCUMULATOR_ADDRESS_TYPE IS STD_LOGIC_VECTOR(ACCUMULATOR_ADDRESS_WIDTH - 1 DOWNTO 0);
    SUBTYPE WEIGHT_ADDRESS_TYPE IS STD_LOGIC_VECTOR(WEIGHT_ADDRESS_WIDTH - 1 DOWNTO 0);
    SUBTYPE LENGTH_TYPE IS STD_LOGIC_VECTOR(LENGTH_WIDTH - 1 DOWNTO 0);
    SUBTYPE OP_CODE_TYPE IS STD_LOGIC_VECTOR(OP_CODE_WIDTH - 1 DOWNTO 0);

    TYPE INSTRUCTION_TYPE IS RECORD
        OP_CODE : OP_CODE_TYPE;
        CALC_LENGTH : LENGTH_TYPE;
        ACC_ADDRESS : ACCUMULATOR_ADDRESS_TYPE;
        BUFFER_ADDRESS : BUFFER_ADDRESS_TYPE;
    END RECORD INSTRUCTION_TYPE;

    TYPE WEIGHT_INSTRUCTION_TYPE IS RECORD
        OP_CODE : OP_CODE_TYPE;
        CALC_LENGTH : LENGTH_TYPE;
        WEIGHT_ADDRESS : WEIGHT_ADDRESS_TYPE;
    END RECORD WEIGHT_INSTRUCTION_TYPE;

    FUNCTION TO_WEIGHT_INSTRUCTION(INSTRUCTION : INSTRUCTION_TYPE) RETURN WEIGHT_INSTRUCTION_TYPE;

    FUNCTION INSTRUCTION_TO_BITS(INSTRUCTION : INSTRUCTION_TYPE) RETURN STD_LOGIC_VECTOR;

    FUNCTION BITS_TO_INSTRUCTION(BITVECTOR : STD_LOGIC_VECTOR(10 * BYTE_WIDTH - 1 DOWNTO 0)) RETURN INSTRUCTION_TYPE;

    FUNCTION INIT_INSTRUCTION RETURN INSTRUCTION_TYPE;
END TPU_PACK;

PACKAGE BODY TPU_PACK IS
    FUNCTION BITS_TO_ACTIVATION(BITVECTOR : ACTIVATION_BIT_TYPE) RETURN ACTIVATION_TYPE IS
    BEGIN
        CASE BITVECTOR IS
            WHEN "0000" => RETURN NO_ACTIVATION;
            WHEN "0001" => RETURN RELU;
            WHEN "0010" => RETURN RELU6;
            WHEN "0011" => RETURN CRELU;
            WHEN "0100" => RETURN ELU;
            WHEN "0101" => RETURN SELU;
            WHEN "0110" => RETURN SOFTPLUS;
            WHEN "0111" => RETURN SOFTSIGN;
            WHEN "1000" => RETURN DROPOUT;
            WHEN "1001" => RETURN SIGMOID;
            WHEN "1010" => RETURN TANH;
            WHEN OTHERS =>
                REPORT "Unknown activation function!" SEVERITY ERROR;
                RETURN NO_ACTIVATION;
        END CASE;
    END FUNCTION BITS_TO_ACTIVATION;

    FUNCTION ACTIVATION_TO_BITS(ACTIVATION_FUNCTION : ACTIVATION_TYPE) RETURN ACTIVATION_BIT_TYPE IS
    BEGIN
        CASE ACTIVATION_FUNCTION IS
            WHEN NO_ACTIVATION => RETURN "0000";
            WHEN RELU => RETURN "0001";
            WHEN RELU6 => RETURN "0010";
            WHEN CRELU => RETURN "0011";
            WHEN ELU => RETURN "0100";
            WHEN SELU => RETURN "0101";
            WHEN SOFTPLUS => RETURN "0110";
            WHEN SOFTSIGN => RETURN "0111";
            WHEN DROPOUT => RETURN "1000";
            WHEN SIGMOID => RETURN "1001";
            WHEN TANH => RETURN "1010";
        END CASE;
    END FUNCTION ACTIVATION_TO_BITS;

    FUNCTION BITS_TO_BYTE_ARRAY(BITVECTOR : STD_LOGIC_VECTOR) RETURN BYTE_ARRAY_TYPE IS
        VARIABLE BYTE_ARRAY : BYTE_ARRAY_TYPE(0 TO ((BITVECTOR'LENGTH / BYTE_WIDTH) - 1));
    BEGIN
        FOR i IN BYTE_ARRAY'RANGE LOOP
            BYTE_ARRAY(i) := BITVECTOR(i * BYTE_WIDTH + BYTE_WIDTH - 1 DOWNTO i * BYTE_WIDTH);
        END LOOP;

        RETURN BYTE_ARRAY;
    END FUNCTION BITS_TO_BYTE_ARRAY;

    FUNCTION BYTE_ARRAY_TO_BITS(BYTE_ARRAY : BYTE_ARRAY_TYPE) RETURN STD_LOGIC_VECTOR IS
        VARIABLE BITVECTOR : STD_LOGIC_VECTOR(((BYTE_ARRAY'LENGTH * BYTE_WIDTH) - 1) DOWNTO 0);
    BEGIN
        FOR i IN BYTE_ARRAY'RANGE LOOP
            BITVECTOR(i * BYTE_WIDTH + BYTE_WIDTH - 1 DOWNTO i * BYTE_WIDTH) := BYTE_ARRAY(i);
        END LOOP;

        RETURN BITVECTOR;
    END FUNCTION BYTE_ARRAY_TO_BITS;

    FUNCTION BITS_TO_WORD_ARRAY(BITVECTOR : STD_LOGIC_VECTOR) RETURN WORD_ARRAY_TYPE IS
        VARIABLE WORD_ARRAY : WORD_ARRAY_TYPE(0 TO ((BITVECTOR'LENGTH / (4 * BYTE_WIDTH)) - 1));
    BEGIN
        FOR i IN WORD_ARRAY'RANGE LOOP
            WORD_ARRAY(i) := BITVECTOR(i * 4 * BYTE_WIDTH + 4 * BYTE_WIDTH - 1 DOWNTO i * 4 * BYTE_WIDTH);
        END LOOP;

        RETURN WORD_ARRAY;
    END FUNCTION BITS_TO_WORD_ARRAY;

    FUNCTION WORD_ARRAY_TO_BITS(WORD_ARRAY : WORD_ARRAY_TYPE) RETURN STD_LOGIC_VECTOR IS
        VARIABLE BITVECTOR : STD_LOGIC_VECTOR(((WORD_ARRAY'LENGTH * 4 * BYTE_WIDTH) - 1) DOWNTO 0);
    BEGIN
        FOR i IN WORD_ARRAY'RANGE LOOP
            BITVECTOR(i * 4 * BYTE_WIDTH + 4 * BYTE_WIDTH - 1 DOWNTO i * 4 * BYTE_WIDTH) := WORD_ARRAY(i);
        END LOOP;

        RETURN BITVECTOR;
    END FUNCTION WORD_ARRAY_TO_BITS;

    FUNCTION TO_WEIGHT_INSTRUCTION(INSTRUCTION : INSTRUCTION_TYPE) RETURN WEIGHT_INSTRUCTION_TYPE IS
        VARIABLE WEIGHT_INSTRUCTION : WEIGHT_INSTRUCTION_TYPE;
    BEGIN
        WEIGHT_INSTRUCTION.OP_CODE := INSTRUCTION.OP_CODE;
        WEIGHT_INSTRUCTION.CALC_LENGTH := INSTRUCTION.CALC_LENGTH;
        WEIGHT_INSTRUCTION.WEIGHT_ADDRESS := INSTRUCTION.BUFFER_ADDRESS & INSTRUCTION.ACC_ADDRESS;

        RETURN WEIGHT_INSTRUCTION;
    END FUNCTION TO_WEIGHT_INSTRUCTION;

    FUNCTION INSTRUCTION_TO_BITS(INSTRUCTION : INSTRUCTION_TYPE) RETURN STD_LOGIC_VECTOR IS
        VARIABLE BITVECTOR : STD_LOGIC_VECTOR(10 * BYTE_WIDTH - 1 DOWNTO 0);
    BEGIN
        BITVECTOR(OP_CODE_WIDTH - 1 DOWNTO 0) := INSTRUCTION.OP_CODE;
        BITVECTOR(LENGTH_WIDTH + OP_CODE_WIDTH - 1 DOWNTO OP_CODE_WIDTH) := INSTRUCTION.CALC_LENGTH;
        BITVECTOR(ACCUMULATOR_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH - 1 DOWNTO LENGTH_WIDTH + OP_CODE_WIDTH) := INSTRUCTION.ACC_ADDRESS;
        BITVECTOR(BUFFER_ADDRESS_WIDTH + ACCUMULATOR_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH - 1 DOWNTO ACCUMULATOR_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH) := INSTRUCTION.BUFFER_ADDRESS;

        RETURN BITVECTOR;
    END FUNCTION INSTRUCTION_TO_BITS;

    FUNCTION BITS_TO_INSTRUCTION(BITVECTOR : STD_LOGIC_VECTOR(10 * BYTE_WIDTH - 1 DOWNTO 0)) RETURN INSTRUCTION_TYPE IS
        VARIABLE INSTRUCTION : INSTRUCTION_TYPE;
    BEGIN
        INSTRUCTION.OP_CODE := BITVECTOR(OP_CODE_WIDTH - 1 DOWNTO 0);
        INSTRUCTION.CALC_LENGTH := BITVECTOR(LENGTH_WIDTH + OP_CODE_WIDTH - 1 DOWNTO OP_CODE_WIDTH);
        INSTRUCTION.ACC_ADDRESS := BITVECTOR(ACCUMULATOR_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH - 1 DOWNTO LENGTH_WIDTH + OP_CODE_WIDTH);
        INSTRUCTION.BUFFER_ADDRESS := BITVECTOR(BUFFER_ADDRESS_WIDTH + ACCUMULATOR_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH - 1 DOWNTO ACCUMULATOR_ADDRESS_WIDTH + LENGTH_WIDTH + OP_CODE_WIDTH);

        RETURN INSTRUCTION;
    END FUNCTION BITS_TO_INSTRUCTION;

    FUNCTION INIT_INSTRUCTION RETURN INSTRUCTION_TYPE IS
    BEGIN
        RETURN (
        OP_CODE => (OTHERS => '0'),
        CALC_LENGTH => (OTHERS => '0'),
        ACC_ADDRESS => (OTHERS => '0'),
        BUFFER_ADDRESS => (OTHERS => '0')
        );
    END FUNCTION INIT_INSTRUCTION;
END PACKAGE BODY;